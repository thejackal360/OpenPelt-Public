.title TEC Model

.INC "output/params.mod"

* TEC thermal resistance. Units: ?
* TODO: TEMP DEPENDENT
.PARAM R_TEC = (L_TEC/(k_TEC^A_TEC))
.PARAM CAP_TEC = (m_TEC^c_TEC)
.PARAM CAP_METAL = (m_METAL^c_METAL)
.PARAM R_METAL = (L_METAL/(k_METAL^A_METAL))

*** Electrical Circuit ***

* Source voltage
a1 %v([tecplus]) filesrc

* Rs - source resistance
R1 tecplus seebeck {Rs}

* Seebeck effect
B1 seebeck tecminus V={alpha}^(v(th)-v(tc))

*** Thermal Circuit ***

* TEC thermal resistance. Units: ?
R2 tc th {R_TEC}

* TEC thermal capacitance. Units: ?
C1 tc th {CAP_TEC}

* Metal thermal capacitance. Units: ?
C2 tamb th {CAP_METAL}

* Metal thermal resistance. Units: ?
R3 tamb th {R_METAL}

* Q_pc heat pumping current. Units: ?
B2 tc tamb I={alpha}^i(R1)^v(tc)

* Ohmic heat current to coldside
B3 tamb tc I=i(R1)^i(R1)^{Rs}/2

* Ohmic heat current to hotside
B4 tamb th I=i(R1)^i(R1)^{Rs}/2

* Q_ph heat pumping current. Units: ?
B5 tamb th I={alpha}^i(R1)^v(th)

*** Control ***
.control
    save v(th)
    tran 10u 10m
    wrdata output v(th)
.endc

.end
