***************************************
* SIMULATION OF MEASURING SYSTEM
* TAMB = AMBIENT TEMPERATURE
* SE = SEEBECK CONSTANT
***************************************
.PARAM TAMB=296.4, SE=0.05292, RM=1.806, RP=1.8
*********************************
******** THERMAL CIRCUIT ********
*********************************
*** HEAT SINK ***
V1 3 0 DC {TAMB}
R1 4 3 0.34
C1 4 0 340 IC={TAMB}
R2 4 1 0.143
*** THERMAL PELTIER MODEL ***
C2 1 0 2 IC={TAMB}
G1 0 1 VALUE={((V(13) - V(12))/{RP})*(((V(13) - V(12))/{RP})*RP+SE*(V(1)-V(2)))}
R3 1 2 1.768
G2 2 1 VALUE={((V(13) - V(12))/{RP})*(SE*V(2)-0.9*((V(13) - V(12))/{RP}))}
C3 2 0 2 IC={TAMB}
*** THERMAL MASS ***
R4 5 2 0.143
C4 5 0 304 IC={TAMB}
R5 5 3 3.1
************************************
******** ELECTRICAL CIRCUIT ********
************************************
*** ELECTRICAL PELTIER MODEL ***
V2 11 13 DC 0
R6 13 12 {RP}
E1 12 0 VALUE = {{SE}*(V(1)-V(2))}
***** EXTERNAL CURRENT SOURCE *****
I1 0 11 2.1
.OPTIONS RELTOL=5U
.CONTROL
    TRAN 1 2K UIC
    SAVE v(2) v(1)
    WRDATA OUTPUT_C v(2)
    WRDATA OUTPUT_H v(1)
    EXIT
.ENDC
.END
*****************************************
